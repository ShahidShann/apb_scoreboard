//write scoreboard check for apb protocol, consider single master and single slave .

class scoreboard extends uvm_scoreboard
  //factory registration
  //declaration of ports from monitor/refrennce model
  //constructor
  //build phase
  //connect phase
  //run phase 
  //write scoreboard check here with expected and actual data
endclass
