class scoreboard extends uvm_scoreboard
  //factory registration
  //declaration of analysis_imp_ports from monitor/refrennce model
  //constructor
  //build phase
  //connect phase
  //run phase 
  //write scorebrd check here with expected and actual data
endclass
